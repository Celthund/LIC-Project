-- TestBench Template 

  LIBRARY ieee;
  USE ieee.std_logic_1164.ALL;
  USE ieee.numeric_std.ALL;

  ENTITY KS_TEST IS
  END KS_TEST;

  ARCHITECTURE behavior OF KS_TEST IS 

  -- Component Declaration
          COMPONENT KeyScan
          PORT( 
					RST: in STD_LOGIC;
					CLK : in  STD_LOGIC;
					KScan : in  STD_LOGIC_VECTOR (1 downto 0);
					K : out  STD_LOGIC_VECTOR (3 downto 0);
					PENC_IN: in  STD_LOGIC_VECTOR (3 downto 0);
					KPress : out  STD_LOGIC;
					DEC_OUT : buffer STD_LOGIC_VECTOR (2 downto 0)
          );
          END COMPONENT;
				
			 -- Inputs
          SIGNAL CLK :  std_logic := '0';
			 SIGNAL RST :  std_logic := '0';
          SIGNAL KScan :  std_logic_vector(1 downto 0);
			 SIGNAL PENC_IN :  std_logic_vector(3 downto 0);
          
			 -- Outputs
			 SIGNAL KPress :  std_logic := '0';
			 SIGNAL DEC_OUT : STD_LOGIC_VECTOR (2 downto 0);
			 SIGNAL K : STD_LOGIC_VECTOR (3 downto 0);
			 
			 -- Clock period definitions
			 constant CLK_period : time := 10 ns;
  BEGIN

  -- Component Instantiation
          uud:  KeyScan PORT MAP(
					RST => RST,
					CLK => CLK,
					KScan => KScan,
					K => K,
					PENC_IN => PENC_IN,
					KPress => KPress,
					DEC_OUT => DEC_OUT
          );

		CLK_process :process
	   begin
			CLK <= '0';
			wait for CLK_period/2;
			CLK <= '1';
			wait for CLK_period/2;
		end process;
	  
  --  Test Bench Statements
     tb : PROCESS
     BEGIN
			RST <= '1';
			KScan <= "00";
			PENC_IN <= "1111";
         wait for 100 ns; -- wait until global set/reset completes
			RST <= '0';
        -- Add user defined stimulus here
			
			-- Test for key presses in first column
			PENC_IN <= "1110";
			
			KScan <= "01";
			wait for CLK_period * 10; -- K <= "0000"; KPress <= '1'
			
			PENC_IN <= "1111";
			KScan <= "00";
			wait for CLK_period * 10; -- Reset; Kpress <= '0'
			
			PENC_IN <= "1101";
			wait for CLK_period;
			KScan <= "01";
			wait for CLK_period * 10; -- K <= "0001"
			
			PENC_IN <= "1111";
			KScan <= "10";
			wait for CLK_period * 10; -- Reset; Kpress <= '0'
			
			-- Test for key presses in first column
			PENC_IN <= "1110";
			KScan <= "01";
			wait for CLK_period * 10; -- K <= "0000"; KPress <= '1'
			
			PENC_IN <= "1111";
			KScan <= "00";
			wait for CLK_period * 10; -- Reset; Kpress <= '0'
			
			
			wait; -- will wait forever
     END PROCESS tb;
  --  End Test Bench 

  END;
